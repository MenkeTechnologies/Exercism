module main

fn truncate(s string) string {
	return s.limit(5)
}

